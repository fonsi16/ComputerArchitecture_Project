`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:06:52 02/29/2024 
// Design Name: 
// Module Name:    Mux_R 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Mux_R(
    input [7:0] Constante,
    input [7:0] Dados_M,
    input [7:0] Dados_IN,
    input [7:0] Resultado,
    output [7:0] Dados_R,
    input [2:0] SEL_Dados
    );


endmodule
